

module round_robin_test